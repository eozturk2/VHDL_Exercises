-- Code your testbench here
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity testbench is
end testbench;

architecture tb of testbench is

component FP_Adder is
port(
	 A,B	: in std_logic_vector(31 downto 0);
     S		: out std_logic_vector(31 downto 0));
end component;

signal A,B	: std_logic_vector(31 downto 0);
signal S	: std_logic_vector(31 downto 0);

-- Test Cases:

-- Sign Test:

-- A = 100.35  = 01000010110010001011001100110011
-- B = 25.58   = 01000001110011001010001111010111
-- S = 125.93  = 01000010111110111101110000101001
-- Actual	     = 01000010111110111101110000101000

-- A = -100.35 = 11000010110010001011001100110011
-- B = 25.58   = 01000001110011001010001111010111
-- S = -74.77  = 11000010100101011000101000111101
-- Actual	     = 11000010100101011000101000111101

-- A = 100.35  = 01000010110010001011001100110011
-- B = -25.58  = 11000001110011001010001111010111
-- S = 74.77   = 01000010100101011000101000111101
-- Actual      = 01000010100101011000101000111101

-- A = -100.35 = 11000010110010001011001100110011
-- B = -25.58  = 11000001110011001010001111010111
-- S = -125.93 = 11000010111110111101110000101001
-- Actual      = 11000010111110111101110000101000

-- Random Large Numbers:

-- A = 18752046.45 = 01001011100011110001000100010111
-- B = 64041767.91 = 01001100011101000100110011001010
-- S = 82793814.36 = 01001100100111011110101010101011
-- Actual          = 01001100100111011110101010101011

-- A = 302369641.84 = 01001101100100000010111001011011
-- B = 45824505.98  = 01001100001011101100111001111110
-- S = 348194147.82 = 01001101101001100000100000101011
-- Actual			      = 01001101101001100000100000101011

-- Special Cases:

-- A = Infinity  = 01111111100000000000000000000000
-- B = Infinity  = 01111111100000000000000000000000
-- S = Infinity  = 01111111100000000000000000000000
-- Actual        = 01111111100000000000000000000000

-- A = -Infinity = 11111111100000000000000000000000
-- B = -Infinity = 11111111100000000000000000000000
-- S = -Infinity = 11111111100000000000000000000000
-- Actual        = 11111111100000000000000000000000

-- A = Infinity  = 01111111100000000000000000000000
-- B = -Infinity = 11111111100000000000000000000000
-- S = NaN		   = 011111111 + (nonzero mantissa)
-- Actual		     = 01111111100000000000000000000001

-- (Same for -inf)
-- A = Infinity  = 01111111100000000000000000000000
-- B = 100.35    = 01000010110010001011001100110011
-- S = Infinity  = 01111111100000000000000000000000
-- Actual		     = 01111111100000000000000000000000
