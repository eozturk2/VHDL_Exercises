-- Code your testbench here
library IEEE;
use IEEE.std_logic_1164.all;

entity testbench is

end testbench;

architecture tb of testbench is

component my_NAND_gate is
port(
	a: in std_logic;
    b: in std_logic;
    q: out std_logic);
end component;

signal a_in, b_in, q_out: std_logic;

begin
	DUT: my_NAND_gate port map (a_in, b_in, q_out);
    process
    begin
    	a_in <= '0';
        b_in <= '0';
        wait for 1 ns;
        
        a_in <= '0';
        b_in <= '1';
        wait for 1 ns;
        
        a_in <= '1';
        b_in <= '0';
        wait for 1 ns;
        
        a_in <= '1';
        b_in <= '1';
        wait for 1 ns;
        
        a_in <= '0';
        b_in <= '0';
        
        wait;
    end process;
end tb;
